module cir
(
    input   a;
    output  b;
    wire    c;
);
    assign 
endmodule